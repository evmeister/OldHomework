library verilog;
use verilog.vl_types.all;
entity parta_vlg_vec_tst is
end parta_vlg_vec_tst;

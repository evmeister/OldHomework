library verilog;
use verilog.vl_types.all;
entity Bigmux_vlg_vec_tst is
end Bigmux_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity parta_vlg_check_tst is
    port(
        LED0            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end parta_vlg_check_tst;

library verilog;
use verilog.vl_types.all;
entity Lab05_vlg_vec_tst is
end Lab05_vlg_vec_tst;

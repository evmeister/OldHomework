`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Evan Eberhardt
// James Olwell
// 
// Create Date: 06/05/2017 05:45:26 PM
// Module Name: CPU
// Project Name: Final Project
//////////////////////////////////////////////////////////////////////////////////


module CPU(

    );
endmodule

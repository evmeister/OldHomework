library verilog;
use verilog.vl_types.all;
entity Lab05_vlg_check_tst is
    port(
        \Out\           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Lab05_vlg_check_tst;
